library verilog;
use verilog.vl_types.all;
entity div_clk_vlg_vec_tst is
end div_clk_vlg_vec_tst;
